library verilog;
use verilog.vl_types.all;
entity MIPS_Multiciclo_vlg_vec_tst is
end MIPS_Multiciclo_vlg_vec_tst;
